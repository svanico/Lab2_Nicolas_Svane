-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Nov 22 14:37:32 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY sec_luces IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        luz1 : OUT STD_LOGIC;
        luz2 : OUT STD_LOGIC;
        luz3 : OUT STD_LOGIC;
        luz4 : OUT STD_LOGIC
    );
END sec_luces;

ARCHITECTURE BEHAVIOR OF sec_luces IS
    TYPE type_fstate IS (state1,state2,state3,state5,state6,state7,state4);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            luz1 <= '0';
            luz2 <= '0';
            luz3 <= '0';
            luz4 <= '0';
        ELSE
            luz1 <= '0';
            luz2 <= '0';
            luz3 <= '0';
            luz4 <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= state2;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    luz3 <= '1';

                    luz1 <= '1';

                    luz2 <= '1';

                    luz4 <= '1';
                WHEN state2 =>
                    reg_fstate <= state3;

                    luz3 <= '0';

                    luz1 <= '1';

                    luz2 <= '0';

                    luz4 <= '1';
                WHEN state3 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= state4;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    luz3 <= '0';

                    luz1 <= '0';

                    luz2 <= '0';

                    luz4 <= '0';
                WHEN state5 =>
                    reg_fstate <= state6;

                    luz3 <= '1';

                    luz1 <= '0';

                    luz2 <= '1';

                    luz4 <= '1';
                WHEN state6 =>
                    reg_fstate <= state3;

                    luz3 <= '1';

                    luz1 <= '0';

                    luz2 <= '1';

                    luz4 <= '0';
                WHEN state7 =>
                    reg_fstate <= state1;

                    luz3 <= '0';

                    luz1 <= '0';

                    luz2 <= '0';

                    luz4 <= '1';
                WHEN state4 =>
                    reg_fstate <= state1;

                    luz3 <= '1';

                    luz1 <= '0';

                    luz2 <= '1';

                    luz4 <= '0';
                WHEN OTHERS => 
                    luz1 <= 'X';
                    luz2 <= 'X';
                    luz3 <= 'X';
                    luz4 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
