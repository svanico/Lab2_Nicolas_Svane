library verilog;
use verilog.vl_types.all;
entity Esquematico_C_vlg_vec_tst is
end Esquematico_C_vlg_vec_tst;
